.title 1.1.2.2
.probe alli

I0 0 out dc 5mA
Ri out 0 {1/2.5m}
R out 0 {1/(5e-4*(4-V(out)))}

.control
op
print all
let U_A = V(out)
let I_A = I(R)
print U_A, I_A
.endc
.end